----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.11.2023 11:20:49
-- Design Name: 
-- Module Name: Init_VGA - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Init_VGA is
    Port ( clk : in STD_LOGIC;
            reset : in STD_LOGIC;
            init_vga : in std_logic;
           write : out std_logic;
           data : out std_logic_vector ( 11 downto 0);
           row : out STD_LOGIC_VECTOR (8 downto 0);
           collumn : out STD_LOGIC_VECTOR (7 downto 0);
           init_complete: out std_logic);
end Init_VGA;

architecture Behavioral of Init_VGA is

TYPE vga_init IS ARRAY (0 TO 3361) OF integer;
signal init: vga_init:= (16, 73, 16, 74, 16, 75, 16, 76, 16, 77, 16, 78, 16, 79, 16, 80, 16, 81, 16, 82, 16, 83, 16, 84, 16, 89, 16, 90, 16, 91, 16, 92, 16, 101, 16, 102, 16, 103, 16, 104, 16, 113, 16, 114, 16, 115, 16, 116, 16, 117, 16, 118, 16, 119, 16, 120, 16, 129, 16, 130, 16, 131, 16, 132, 16, 141, 16, 142, 16, 143, 16, 144, 16, 149, 16, 150, 16, 151, 16, 152, 16, 153, 16, 154, 16, 155, 16, 156, 16, 157, 16, 158, 16, 159, 16, 160, 16, 161, 16, 162, 16, 163, 16, 164, 16, 181, 16, 182, 16, 183, 16, 184, 16, 185, 16, 186, 16, 187, 16, 188, 16, 201, 16, 202, 16, 203, 16, 204, 16, 205, 16, 206, 16, 207, 16, 208, 16, 217, 16, 218, 16, 219, 16, 220, 16, 233, 16, 234, 16, 235, 16, 236, 16, 241, 16, 242, 16, 243, 16, 244, 16, 245, 16, 246, 16, 247, 16, 248, 16, 249, 16, 250, 16, 251, 16, 252, 16, 253, 16, 254, 16, 255, 16, 256, 17, 73, 17, 74, 17, 75, 17, 76, 17, 77, 17, 78, 17, 79, 17, 80, 17, 81, 17, 82, 17, 83, 17, 84, 17, 89, 17, 90, 17, 91, 17, 92, 17, 101, 17, 102, 17, 103, 17, 104, 17, 113, 17, 114, 17, 115, 17, 116, 17, 117, 17, 118, 17, 119, 17, 120, 17, 129, 17, 130, 17, 131, 17, 132, 17, 141, 17, 142, 17, 143, 17, 144, 17, 149, 17, 150, 17, 151, 17, 152, 17, 153, 17, 154, 17, 155, 17, 156, 17, 157, 17, 158, 17, 159, 17, 160, 17, 161, 17, 162, 17, 163, 17, 164, 17, 181, 17, 182, 17, 183, 17, 184, 17, 185, 17, 186, 17, 187, 17, 188, 17, 201, 17, 202, 17, 203, 17, 204, 17, 205, 17, 206, 17, 207, 17, 208, 17, 217, 17, 218, 17, 219, 17, 220, 17, 233, 17, 234, 17, 235, 17, 236, 17, 241, 17, 242, 17, 243, 17, 244, 17, 245, 17, 246, 17, 247, 17, 248, 17, 249, 17, 250, 17, 251, 17, 252, 17, 253, 17, 254, 17, 255, 17, 256, 18, 73, 18, 74, 18, 75, 18, 76, 18, 77, 18, 78, 18, 79, 18, 80, 18, 81, 18, 82, 18, 83, 18, 84, 18, 89, 18, 90, 18, 91, 18, 92, 18, 101, 18, 102, 18, 103, 18, 104, 18, 113, 18, 114, 18, 115, 18, 116, 18, 117, 18, 118, 18, 119, 18, 120, 18, 129, 18, 130, 18, 131, 18, 132, 18, 141, 18, 142, 18, 143, 18, 144, 18, 149, 18, 150, 18, 151, 18, 152, 18, 153, 18, 154, 18, 155, 18, 156, 18, 157, 18, 158, 18, 159, 18, 160, 18, 161, 18, 162, 18, 163, 18, 164, 18, 181, 18, 182, 18, 183, 18, 184, 18, 185, 18, 186, 18, 187, 18, 188, 18, 201, 18, 202, 18, 203, 18, 204, 18, 205, 18, 206, 18, 207, 18, 208, 18, 217, 18, 218, 18, 219, 18, 220, 18, 233, 18, 234, 18, 235, 18, 236, 18, 241, 18, 242, 18, 243, 18, 244, 18, 245, 18, 246, 18, 247, 18, 248, 18, 249, 18, 250, 18, 251, 18, 252, 18, 253, 18, 254, 18, 255, 18, 256, 19, 73, 19, 74, 19, 75, 19, 76, 19, 77, 19, 78, 19, 79, 19, 80, 19, 81, 19, 82, 19, 83, 19, 84, 19, 89, 19, 90, 19, 91, 19, 92, 19, 101, 19, 102, 19, 103, 19, 104, 19, 113, 19, 114, 19, 115, 19, 116, 19, 117, 19, 118, 19, 119, 19, 120, 19, 129, 19, 130, 19, 131, 19, 132, 19, 141, 19, 142, 19, 143, 19, 144, 19, 149, 19, 150, 19, 151, 19, 152, 19, 153, 19, 154, 19, 155, 19, 156, 19, 157, 19, 158, 19, 159, 19, 160, 19, 161, 19, 162, 19, 163, 19, 164, 19, 181, 19, 182, 19, 183, 19, 184, 19, 185, 19, 186, 19, 187, 19, 188, 19, 201, 19, 202, 19, 203, 19, 204, 19, 205, 19, 206, 19, 207, 19, 208, 19, 217, 19, 218, 19, 219, 19, 220, 19, 233, 19, 234, 19, 235, 19, 236, 19, 241, 19, 242, 19, 243, 19, 244, 19, 245, 19, 246, 19, 247, 19, 248, 19, 249, 19, 250, 19, 251, 19, 252, 19, 253, 19, 254, 19, 255, 19, 256, 20, 69, 20, 70, 20, 71, 20, 72, 20, 89, 20, 90, 20, 91, 20, 92, 20, 93, 20, 94, 20, 95, 20, 96, 20, 101, 20, 102, 20, 103, 20, 104, 20, 109, 20, 110, 20, 111, 20, 112, 20, 121, 20, 122, 20, 123, 20, 124, 20, 129, 20, 130, 20, 131, 20, 132, 20, 137, 20, 138, 20, 139, 20, 140, 20, 149, 20, 150, 20, 151, 20, 152, 20, 177, 20, 178, 20, 179, 20, 180, 20, 197, 20, 198, 20, 199, 20, 200, 20, 209, 20, 210, 20, 211, 20, 212, 20, 217, 20, 218, 20, 219, 20, 220, 20, 221, 20, 222, 20, 223, 20, 224, 20, 229, 20, 230, 20, 231, 20, 232, 20, 233, 20, 234, 20, 235, 20, 236, 20, 241, 20, 242, 20, 243, 20, 244, 21, 69, 21, 70, 21, 71, 21, 72, 21, 89, 21, 90, 21, 91, 21, 92, 21, 93, 21, 94, 21, 95, 21, 96, 21, 101, 21, 102, 21, 103, 21, 104, 21, 109, 21, 110, 21, 111, 21, 112, 21, 121, 21, 122, 21, 123, 21, 124, 21, 129, 21, 130, 21, 131, 21, 132, 21, 137, 21, 138, 21, 139, 21, 140, 21, 149, 21, 150, 21, 151, 21, 152, 21, 177, 21, 178, 21, 179, 21, 180, 21, 197, 21, 198, 21, 199, 21, 200, 21, 209, 21, 210, 21, 211, 21, 212, 21, 217, 21, 218, 21, 219, 21, 220, 21, 221, 21, 222, 21, 223, 21, 224, 21, 229, 21, 230, 21, 231, 21, 232, 21, 233, 21, 234, 21, 235, 21, 236, 21, 241, 21, 242, 21, 243, 21, 244, 22, 69, 22, 70, 22, 71, 22, 72, 22, 89, 22, 90, 22, 91, 22, 92, 22, 93, 22, 94, 22, 95, 22, 96, 22, 101, 22, 102, 22, 103, 22, 104, 22, 109, 22, 110, 22, 111, 22, 112, 22, 121, 22, 122, 22, 123, 22, 124, 22, 129, 22, 130, 22, 131, 22, 132, 22, 137, 22, 138, 22, 139, 22, 140, 22, 149, 22, 150, 22, 151, 22, 152, 22, 177, 22, 178, 22, 179, 22, 180, 22, 197, 22, 198, 22, 199, 22, 200, 22, 209, 22, 210, 22, 211, 22, 212, 22, 217, 22, 218, 22, 219, 22, 220, 22, 221, 22, 222, 22, 223, 22, 224, 22, 229, 22, 230, 22, 231, 22, 232, 22, 233, 22, 234, 22, 235, 22, 236, 22, 241, 22, 242, 22, 243, 22, 244, 23, 69, 23, 70, 23, 71, 23, 72, 23, 89, 23, 90, 23, 91, 23, 92, 23, 93, 23, 94, 23, 95, 23, 96, 23, 101, 23, 102, 23, 103, 23, 104, 23, 109, 23, 110, 23, 111, 23, 112, 23, 121, 23, 122, 23, 123, 23, 124, 23, 129, 23, 130, 23, 131, 23, 132, 23, 137, 23, 138, 23, 139, 23, 140, 23, 149, 23, 150, 23, 151, 23, 152, 23, 177, 23, 178, 23, 179, 23, 180, 23, 197, 23, 198, 23, 199, 23, 200, 23, 209, 23, 210, 23, 211, 23, 212, 23, 217, 23, 218, 23, 219, 23, 220, 23, 221, 23, 222, 23, 223, 23, 224, 23, 229, 23, 230, 23, 231, 23, 232, 23, 233, 23, 234, 23, 235, 23, 236, 23, 241, 23, 242, 23, 243, 23, 244, 24, 73, 24, 74, 24, 75, 24, 76, 24, 77, 24, 78, 24, 79, 24, 80, 24, 89, 24, 90, 24, 91, 24, 92, 24, 97, 24, 98, 24, 99, 24, 100, 24, 101, 24, 102, 24, 103, 24, 104, 24, 109, 24, 110, 24, 111, 24, 112, 24, 113, 24, 114, 24, 115, 24, 116, 24, 117, 24, 118, 24, 119, 24, 120, 24, 121, 24, 122, 24, 123, 24, 124, 24, 129, 24, 130, 24, 131, 24, 132, 24, 133, 24, 134, 24, 135, 24, 136, 24, 149, 24, 150, 24, 151, 24, 152, 24, 153, 24, 154, 24, 155, 24, 156, 24, 157, 24, 158, 24, 159, 24, 160, 24, 177, 24, 178, 24, 179, 24, 180, 24, 185, 24, 186, 24, 187, 24, 188, 24, 189, 24, 190, 24, 191, 24, 192, 24, 197, 24, 198, 24, 199, 24, 200, 24, 201, 24, 202, 24, 203, 24, 204, 24, 205, 24, 206, 24, 207, 24, 208, 24, 209, 24, 210, 24, 211, 24, 212, 24, 217, 24, 218, 24, 219, 24, 220, 24, 225, 24, 226, 24, 227, 24, 228, 24, 233, 24, 234, 24, 235, 24, 236, 24, 241, 24, 242, 24, 243, 24, 244, 24, 245, 24, 246, 24, 247, 24, 248, 24, 249, 24, 250, 24, 251, 24, 252, 25, 73, 25, 74, 25, 75, 25, 76, 25, 77, 25, 78, 25, 79, 25, 80, 25, 89, 25, 90, 25, 91, 25, 92, 25, 97, 25, 98, 25, 99, 25, 100, 25, 101, 25, 102, 25, 103, 25, 104, 25, 109, 25, 110, 25, 111, 25, 112, 25, 113, 25, 114, 25, 115, 25, 116, 25, 117, 25, 118, 25, 119, 25, 120, 25, 121, 25, 122, 25, 123, 25, 124, 25, 129, 25, 130, 25, 131, 25, 132, 25, 133, 25, 134, 25, 135, 25, 136, 25, 149, 25, 150, 25, 151, 25, 152, 25, 153, 25, 154, 25, 155, 25, 156, 25, 157, 25, 158, 25, 159, 25, 160, 25, 177, 25, 178, 25, 179, 25, 180, 25, 185, 25, 186, 25, 187, 25, 188, 25, 189, 25, 190, 25, 191, 25, 192, 25, 197, 25, 198, 25, 199, 25, 200, 25, 201, 25, 202, 25, 203, 25, 204, 25, 205, 25, 206, 25, 207, 25, 208, 25, 209, 25, 210, 25, 211, 25, 212, 25, 217, 25, 218, 25, 219, 25, 220, 25, 225, 25, 226, 25, 227, 25, 228, 25, 233, 25, 234, 25, 235, 25, 236, 25, 241, 25, 242, 25, 243, 25, 244, 25, 245, 25, 246, 25, 247, 25, 248, 25, 249, 25, 250, 25, 251, 25, 252, 26, 73, 26, 74, 26, 75, 26, 76, 26, 77, 26, 78, 26, 79, 26, 80, 26, 89, 26, 90, 26, 91, 26, 92, 26, 97, 26, 98, 26, 99, 26, 100, 26, 101, 26, 102, 26, 103, 26, 104, 26, 109, 26, 110, 26, 111, 26, 112, 26, 113, 26, 114, 26, 115, 26, 116, 26, 117, 26, 118, 26, 119, 26, 120, 26, 121, 26, 122, 26, 123, 26, 124, 26, 129, 26, 130, 26, 131, 26, 132, 26, 133, 26, 134, 26, 135, 26, 136, 26, 149, 26, 150, 26, 151, 26, 152, 26, 153, 26, 154, 26, 155, 26, 156, 26, 157, 26, 158, 26, 159, 26, 160, 26, 177, 26, 178, 26, 179, 26, 180, 26, 185, 26, 186, 26, 187, 26, 188, 26, 189, 26, 190, 26, 191, 26, 192, 26, 197, 26, 198, 26, 199, 26, 200, 26, 201, 26, 202, 26, 203, 26, 204, 26, 205, 26, 206, 26, 207, 26, 208, 26, 209, 26, 210, 26, 211, 26, 212, 26, 217, 26, 218, 26, 219, 26, 220, 26, 225, 26, 226, 26, 227, 26, 228, 26, 233, 26, 234, 26, 235, 26, 236, 26, 241, 26, 242, 26, 243, 26, 244, 26, 245, 26, 246, 26, 247, 26, 248, 26, 249, 26, 250, 26, 251, 26, 252, 27, 73, 27, 74, 27, 75, 27, 76, 27, 77, 27, 78, 27, 79, 27, 80, 27, 89, 27, 90, 27, 91, 27, 92, 27, 97, 27, 98, 27, 99, 27, 100, 27, 101, 27, 102, 27, 103, 27, 104, 27, 109, 27, 110, 27, 111, 27, 112, 27, 113, 27, 114, 27, 115, 27, 116, 27, 117, 27, 118, 27, 119, 27, 120, 27, 121, 27, 122, 27, 123, 27, 124, 27, 129, 27, 130, 27, 131, 27, 132, 27, 133, 27, 134, 27, 135, 27, 136, 27, 149, 27, 150, 27, 151, 27, 152, 27, 153, 27, 154, 27, 155, 27, 156, 27, 157, 27, 158, 27, 159, 27, 160, 27, 177, 27, 178, 27, 179, 27, 180, 27, 185, 27, 186, 27, 187, 27, 188, 27, 189, 27, 190, 27, 191, 27, 192, 27, 197, 27, 198, 27, 199, 27, 200, 27, 201, 27, 202, 27, 203, 27, 204, 27, 205, 27, 206, 27, 207, 27, 208, 27, 209, 27, 210, 27, 211, 27, 212, 27, 217, 27, 218, 27, 219, 27, 220, 27, 225, 27, 226, 27, 227, 27, 228, 27, 233, 27, 234, 27, 235, 27, 236, 27, 241, 27, 242, 27, 243, 27, 244, 27, 245, 27, 246, 27, 247, 27, 248, 27, 249, 27, 250, 27, 251, 27, 252, 28, 81, 28, 82, 28, 83, 28, 84, 28, 89, 28, 90, 28, 91, 28, 92, 28, 101, 28, 102, 28, 103, 28, 104, 28, 109, 28, 110, 28, 111, 28, 112, 28, 121, 28, 122, 28, 123, 28, 124, 28, 129, 28, 130, 28, 131, 28, 132, 28, 137, 28, 138, 28, 139, 28, 140, 28, 149, 28, 150, 28, 151, 28, 152, 28, 177, 28, 178, 28, 179, 28, 180, 28, 189, 28, 190, 28, 191, 28, 192, 28, 197, 28, 198, 28, 199, 28, 200, 28, 209, 28, 210, 28, 211, 28, 212, 28, 217, 28, 218, 28, 219, 28, 220, 28, 233, 28, 234, 28, 235, 28, 236, 28, 241, 28, 242, 28, 243, 28, 244, 29, 81, 29, 82, 29, 83, 29, 84, 29, 89, 29, 90, 29, 91, 29, 92, 29, 101, 29, 102, 29, 103, 29, 104, 29, 109, 29, 110, 29, 111, 29, 112, 29, 121, 29, 122, 29, 123, 29, 124, 29, 129, 29, 130, 29, 131, 29, 132, 29, 137, 29, 138, 29, 139, 29, 140, 29, 149, 29, 150, 29, 151, 29, 152, 29, 177, 29, 178, 29, 179, 29, 180, 29, 189, 29, 190, 29, 191, 29, 192, 29, 197, 29, 198, 29, 199, 29, 200, 29, 209, 29, 210, 29, 211, 29, 212, 29, 217, 29, 218, 29, 219, 29, 220, 29, 233, 29, 234, 29, 235, 29, 236, 29, 241, 29, 242, 29, 243, 29, 244, 30, 81, 30, 82, 30, 83, 30, 84, 30, 89, 30, 90, 30, 91, 30, 92, 30, 101, 30, 102, 30, 103, 30, 104, 30, 109, 30, 110, 30, 111, 30, 112, 30, 121, 30, 122, 30, 123, 30, 124, 30, 129, 30, 130, 30, 131, 30, 132, 30, 137, 30, 138, 30, 139, 30, 140, 30, 149, 30, 150, 30, 151, 30, 152, 30, 177, 30, 178, 30, 179, 30, 180, 30, 189, 30, 190, 30, 191, 30, 192, 30, 197, 30, 198, 30, 199, 30, 200, 30, 209, 30, 210, 30, 211, 30, 212, 30, 217, 30, 218, 30, 219, 30, 220, 30, 233, 30, 234, 30, 235, 30, 236, 30, 241, 30, 242, 30, 243, 30, 244, 31, 81, 31, 82, 31, 83, 31, 84, 31, 89, 31, 90, 31, 91, 31, 92, 31, 101, 31, 102, 31, 103, 31, 104, 31, 109, 31, 110, 31, 111, 31, 112, 31, 121, 31, 122, 31, 123, 31, 124, 31, 129, 31, 130, 31, 131, 31, 132, 31, 137, 31, 138, 31, 139, 31, 140, 31, 149, 31, 150, 31, 151, 31, 152, 31, 177, 31, 178, 31, 179, 31, 180, 31, 189, 31, 190, 31, 191, 31, 192, 31, 197, 31, 198, 31, 199, 31, 200, 31, 209, 31, 210, 31, 211, 31, 212, 31, 217, 31, 218, 31, 219, 31, 220, 31, 233, 31, 234, 31, 235, 31, 236, 31, 241, 31, 242, 31, 243, 31, 244, 32, 69, 32, 70, 32, 71, 32, 72, 32, 73, 32, 74, 32, 75, 32, 76, 32, 77, 32, 78, 32, 79, 32, 80, 32, 89, 32, 90, 32, 91, 32, 92, 32, 101, 32, 102, 32, 103, 32, 104, 32, 109, 32, 110, 32, 111, 32, 112, 32, 121, 32, 122, 32, 123, 32, 124, 32, 129, 32, 130, 32, 131, 32, 132, 32, 141, 32, 142, 32, 143, 32, 144, 32, 149, 32, 150, 32, 151, 32, 152, 32, 153, 32, 154, 32, 155, 32, 156, 32, 157, 32, 158, 32, 159, 32, 160, 32, 161, 32, 162, 32, 163, 32, 164, 32, 181, 32, 182, 32, 183, 32, 184, 32, 185, 32, 186, 32, 187, 32, 188, 32, 197, 32, 198, 32, 199, 32, 200, 32, 209, 32, 210, 32, 211, 32, 212, 32, 217, 32, 218, 32, 219, 32, 220, 32, 233, 32, 234, 32, 235, 32, 236, 32, 241, 32, 242, 32, 243, 32, 244, 32, 245, 32, 246, 32, 247, 32, 248, 32, 249, 32, 250, 32, 251, 32, 252, 32, 253, 32, 254, 32, 255, 32, 256, 33, 69, 33, 70, 33, 71, 33, 72, 33, 73, 33, 74, 33, 75, 33, 76, 33, 77, 33, 78, 33, 79, 33, 80, 33, 89, 33, 90, 33, 91, 33, 92, 33, 101, 33, 102, 33, 103, 33, 104, 33, 109, 33, 110, 33, 111, 33, 112, 33, 121, 33, 122, 33, 123, 33, 124, 33, 129, 33, 130, 33, 131, 33, 132, 33, 141, 33, 142, 33, 143, 33, 144, 33, 149, 33, 150, 33, 151, 33, 152, 33, 153, 33, 154, 33, 155, 33, 156, 33, 157, 33, 158, 33, 159, 33, 160, 33, 161, 33, 162, 33, 163, 33, 164, 33, 181, 33, 182, 33, 183, 33, 184, 33, 185, 33, 186, 33, 187, 33, 188, 33, 197, 33, 198, 33, 199, 33, 200, 33, 209, 33, 210, 33, 211, 33, 212, 33, 217, 33, 218, 33, 219, 33, 220, 33, 233, 33, 234, 33, 235, 33, 236, 33, 241, 33, 242, 33, 243, 33, 244, 33, 245, 33, 246, 33, 247, 33, 248, 33, 249, 33, 250, 33, 251, 33, 252, 33, 253, 33, 254, 33, 255, 33, 256, 34, 69, 34, 70, 34, 71, 34, 72, 34, 73, 34, 74, 34, 75, 34, 76, 34, 77, 34, 78, 34, 79, 34, 80, 34, 89, 34, 90, 34, 91, 34, 92, 34, 101, 34, 102, 34, 103, 34, 104, 34, 109, 34, 110, 34, 111, 34, 112, 34, 121, 34, 122, 34, 123, 34, 124, 34, 129, 34, 130, 34, 131, 34, 132, 34, 141, 34, 142, 34, 143, 34, 144, 34, 149, 34, 150, 34, 151, 34, 152, 34, 153, 34, 154, 34, 155, 34, 156, 34, 157, 34, 158, 34, 159, 34, 160, 34, 161, 34, 162, 34, 163, 34, 164, 34, 181, 34, 182, 34, 183, 34, 184, 34, 185, 34, 186, 34, 187, 34, 188, 34, 197, 34, 198, 34, 199, 34, 200, 34, 209, 34, 210, 34, 211, 34, 212, 34, 217, 34, 218, 34, 219, 34, 220, 34, 233, 34, 234, 34, 235, 34, 236, 34, 241, 34, 242, 34, 243, 34, 244, 34, 245, 34, 246, 34, 247, 34, 248, 34, 249, 34, 250, 34, 251, 34, 252, 34, 253, 34, 254, 34, 255, 34, 256, 35, 69, 35, 70, 35, 71, 35, 72, 35, 73, 35, 74, 35, 75, 35, 76, 35, 77, 35, 78, 35, 79, 35, 80, 35, 89, 35, 90, 35, 91, 35, 92, 35, 101, 35, 102, 35, 103, 35, 104, 35, 109, 35, 110, 35, 111, 35, 112, 35, 121, 35, 122, 35, 123, 35, 124, 35, 129, 35, 130, 35, 131, 35, 132, 35, 141, 35, 142, 35, 143, 35, 144, 35, 149, 35, 150, 35, 151, 35, 152, 35, 153, 35, 154, 35, 155, 35, 156, 35, 157, 35, 158, 35, 159, 35, 160, 35, 161, 35, 162, 35, 163, 35, 164, 35, 181, 35, 182, 35, 183, 35, 184, 35, 185, 35, 186, 35, 187, 35, 188, 35, 197, 35, 198, 35, 199, 35, 200, 35, 209, 35, 210, 35, 211, 35, 212, 35, 217, 35, 218, 35, 219, 35, 220, 35, 233, 35, 234, 35, 235, 35, 236, 35, 241, 35, 242, 35, 243, 35, 244, 35, 245, 35, 246, 35, 247, 35, 248, 35, 249, 35, 250, 35, 251, 35, 252, 35, 253, 35, 254, 35, 255, 35, 256,51,132); 
signal i_cl : integer :=0;
signal x : integer := 2 ;
signal y : integer := 2;
signal s_write : std_logic;
signal s_data : std_logic_vector(11 downto 0);
begin

process(clk,reset,init_vga)
begin
    if (reset ='1' or init_vga='1') then
        i_cl<=0;
        init_complete <='0';
    elsif(clk'event and clk='1') then
        if(i_cl < 33330) then
            i_cl <= i_cl+1;
             s_write <= '1';
             init_complete <='0';
         else
             init_complete <='1';
        end if;
    end if;
end process;


process(clk, reset, i_cl)
begin
   if (clk'event and clk='1') then
     if (reset ='1' or init_vga ='1') then
        x<=0;
        y<=0;
     elsif (i_cl <1681) then
        y<= init(i_cl*2);
        x<= init(i_cl*2+1);
    else
    
        if(x<=230  ) then
            x <= x + 1;
        else 
            x <= 70;
            if (y < 230) then
                y <= y +1;
            else
                y <=70;
             end if;
         end if;
    end if;
    end if;
end process;

process(x,y)
begin
    if (y<36) then
        if (x<86) or ( x<194 and x>175) then
            s_data <= "000011000000"; 
        else 
            s_data <= "111111111111";           
         end if;
    elsif ((y>=70 and x=230 and y<=230) or (y>=70 and x=70 and y<=230)   or (x>=70 and y=230 and x<=230) or (x>=70 and y=70 and x<=230)) then
        s_data <= "000000001111";
    elsif (y=100 and x<120 and x>=115 ) then
        s_data <= "000011110000";
    elsif (x<230 and x>70 and y<230 and y>70) then
        s_data <= "111111111111";
     else
        s_data <= "000000000000";
    end if;
end process;

data <= s_data;
write <= s_write;
row <= std_logic_vector(to_unsigned(x,9));
collumn <= std_logic_vector(to_unsigned(y,8));


end Behavioral;


